`include "NPU.v"
`include "npu_controller.v"
`include "pe_control_weight.v"
`include "pe_control.v"
`include "pe_result_cache.v"
`include "pe_array.v"
`include "pe.v"
`include "ram_rd_control.v"
`include "ram_wr_control.v"
`include "result_ram.v"
`include "dual_port_ram.v"
