`ifndef AGENT_PKG_SVH
`define AGENT_PKG_SVH

`include "npu_transaction.sv"
`include "npu_master_driver.sv"
`include "npu_master_sequencer.sv"
`include "npu_master_agent.sv"

`endif
