`ifndef NPU_SEQ_SVH
`define NPU_SEQ_SVH

`include "npu_virtual_seq.sv"
`include "npu_sequence.sv"

`endif
