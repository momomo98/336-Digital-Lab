
package npu_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "npu_agent.svh"
    `include "npu_virtual_sequencer.sv"
    `include "npu_seq.svh"
    `include "npu_cov.sv"
    `include "npu_env.sv"
    `include "npu_test.svh"



endpackage




