`ifndef NPU_TEST_SVH
`define NPU_TEST_SVH

`include "npu_base_test.sv"
`include "npu_random_test.sv"

`endif
